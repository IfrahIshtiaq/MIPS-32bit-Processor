module register_file(
    input clk,
    input reset,
    input reg_write_en,
    input [4:0] reg_write_dest,
    input [31:0] reg_write_data,
    input [4:0] reg_read_addr_1,
    output [31:0] reg_read_data_1,
    input [4:0] reg_read_addr_2,
    output [31:0] reg_read_data_2
    );
	 
	 reg     [31:0]     regMem [31:0];  
      // write port  
      //reg [2:0] i;
		initial  
			begin
					   regMem[0]  <= 32'b 000000000000000000000000000000;
						regMem[1]  <= 32'b 000000000000000000000000000001;
						regMem[2]  <= 32'b 000000000000000000000000000010;
						regMem[3]  <= 32'b 000000000000000000000000000011;
						regMem[4]  <= 32'b 000000000000000000000000000100;
						regMem[5]  <= 32'b 000000000000000000000000000101;
						regMem[6]  <= 32'b 000000000000000000000000000110;
						regMem[7]  <= 32'b 000000000000000000000000000111;
						regMem[8]  <= 32'b 000000000000000000000000001000;
						regMem[9]  <= 32'b 000000000000000000000000001001;
						regMem[10]  <= 32'b 000000000000000000000000001010;
						regMem[11]  <= 32'b 000000000000000000000000001011;
						regMem[12]  <= 32'b 000000000000000000000000001100;
						regMem[13]  <= 32'b 000000000000000000000000001101;
						regMem[14]  <= 32'b 000000000000000000000000001110;
						regMem[15]  <= 32'b 000000000000000000000000001111;
						regMem[16]  <= 32'b 000000000000000000000000010000;
						regMem[17]  <= 32'b 000000000000000000000000010001;
						regMem[18]  <= 32'b 000000000000000000000000010010;
						regMem[19]  <= 32'b 000000000000000000000000010011;
						regMem[20]  <= 32'b 000000000000000000000000010100;
						regMem[21]  <= 32'b 000000000000000000000000010101;
						regMem[22]  <= 32'b 000000000000000000000000010110;
						regMem[23]  <= 32'b 000000000000000000000000010111;
						regMem[24]  <= 32'b 000000000000000000000000011000;
						regMem[25]  <= 32'b 000000000000000000000000011001;
						regMem[26]  <= 32'b 000000000000000000000000011010;
						regMem[27]  <= 32'b 000000000000000000000000011011;
						regMem[28]  <= 32'b 000000000000000000000000011100;
						regMem[29]  <= 32'b 000000000000000000000000011101;
						regMem[30]  <= 32'b 000000000000000000000000011110;
						regMem[31]  <= 32'b 000000000000000000000000011111;


				end
      /*always @ (posedge clk or posedge reset) 
			begin  
				if(reset) begin
                regMem[0]  <= 32'b00000000000000000000000000000000;
					 regMem[1]  <= 32'b00000000000000000000000000000000;
				    regMem[2]  <= 32'b00000000000000000000000000000000;
				    regMem[3]  <= 32'b00000000000000000000000000000000;
					 regMem[4]  <= 32'b00000000000000000000000000000000;
					 regMem[5]  <= 32'b00000000000000000000000000000000;
					 regMem[6]  <= 32'b00000000000000000000000000000000;
					 regMem[7]  <= 32'b00000000000000000000000000000000;
					 regMem[8]  <= 32'b00000000000000000000000000000000;
					 regMem[9]  <= 32'b00000000000000000000000000000000;
					 regMem[10] <= 32'b00000000000000000000000000000000;
					 regMem[11] <= 32'b00000000000000000000000000000000;
				    regMem[12] <= 32'b00000000000000000000000000000000;
				    regMem[13] <= 32'b00000000000000000000000000000000;
					 regMem[14] <= 32'b00000000000000000000000000000000;
					 regMem[15] <= 32'b00000000000000000000000000000000;
					 regMem[16] <= 32'b00000000000000000000000000000000;
					 regMem[17] <= 32'b00000000000000000000000000000000;
					 regMem[18] <= 32'b00000000000000000000000000000000;
					 regMem[19] <= 32'b00000000000000000000000000000000;
					 regMem[20] <= 32'b00000000000000000000000000000000;
					 regMem[21] <= 32'b00000000000000000000000000000000;
				    regMem[22] <= 32'b00000000000000000000000000000000;
				    regMem[23] <= 32'b00000000000000000000000000000000;
					 regMem[24] <= 32'b00000000000000000000000000000000;
					 regMem[25] <= 32'b00000000000000000000000000000000;
					 regMem[26] <= 32'b00000000000000000000000000000000;
					 regMem[27] <= 32'b00000000000000000000000000000000;
					 regMem[28] <= 32'b00000000000000000000000000000000;
					 regMem[29] <= 32'b00000000000000000000000000000000;
					 regMem[30] <= 32'b00000000000000000000000000000000;
					 regMem[31] <= 32'b00000000000000000000000000000000;
					 
					 end
    
             else 
						begin  
							 if(reg_write_en) begin  
									regMem[reg_write_dest] <= reg_write_data;  
							 end  
						end    
           end*/
        
      assign reg_read_data_1 = ( reg_read_addr_1 == 0)? 32'b0 : regMem[reg_read_addr_1];  
      assign reg_read_data_2 = ( reg_read_addr_2 == 0)? 32'b0 : regMem[reg_read_addr_2];


endmodule